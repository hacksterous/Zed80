//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.02
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Created Time: Tue May  7 11:16:25 2024

module ROM8kB (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [12:0] ad;

wire [29:0] prom_inst_0_dout_w;
wire [29:0] prom_inst_1_dout_w;
wire [29:0] prom_inst_2_dout_w;
wire [29:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[29:0],dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 2;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hC6508E5D4E808E0ED381CE7381CE39746350FFFFFFFFFFFFFFCBFFC3FFCFFF0F;
defparam prom_inst_0.INIT_RAM_01 = 256'hC39309BADBCEE04146182055E4E8EC63814553CE48E5D8F3578E818E4E1B0739;
defparam prom_inst_0.INIT_RAM_02 = 256'hB5B549FE17894D156D7054DBFFFFFF0DCB3024C672C0F92525C26C63B021FEB6;
defparam prom_inst_0.INIT_RAM_03 = 256'h613B4DB5565B6178F597D3A9390B95B55758B9BC6E54D22FE49365AD586DB5A3;
defparam prom_inst_0.INIT_RAM_04 = 256'h52103912041CFDB8C95070D3F0C1B5424BFB518351C0364F9B82637602095A34;
defparam prom_inst_0.INIT_RAM_05 = 256'h0761EC6D01F3D925BDF1F241706B1CCD6A469FDB3699B3C41650494406B89311;
defparam prom_inst_0.INIT_RAM_06 = 256'hE427353521927FC1F0A9FC25AB7926F1AC9B9C4CE9033AC24D99F1CE53342F26;
defparam prom_inst_0.INIT_RAM_07 = 256'h0AE0B15566AA85FC0544068DD49B416AE17E27C7CA1C1C0503609098108FD188;
defparam prom_inst_0.INIT_RAM_08 = 256'hFB000003533E2E113A5736362169012C8C8C938D3A0D9B3CF4130E17BE3EBAFB;
defparam prom_inst_0.INIT_RAM_09 = 256'h68669721728ED2652793FCAD5D34B445D70BE17B86E4135A09F090BA47E60C30;
defparam prom_inst_0.INIT_RAM_0A = 256'h556D565E565564556E46F6D2712B66045B5E46B49E55E679EC1C4AB49A69A492;
defparam prom_inst_0.INIT_RAM_0B = 256'hE4D7BBCEE4397BF5BBFD6BBBE54BFE27BFD379155DE495E46B5FA7B59EA56957;
defparam prom_inst_0.INIT_RAM_0C = 256'h6AE9ACECBDAB98A258ECFE4B9E5E57925BF2814E5E59E574827B39EFFCE1333E;
defparam prom_inst_0.INIT_RAM_0D = 256'h632EEA23AA6BA8ED5DD276E7A66BD5888E6EDEE4E8BAFBE9BA66B9959598A22A;
defparam prom_inst_0.INIT_RAM_0E = 256'hD8B26C98F4ECB91BE4B2C6DBB046D89EF5E7EE77FE6DB6E7A7618B19BB858F2E;
defparam prom_inst_0.INIT_RAM_0F = 256'h59508D07A02CEE8958B291D6FB9D23F2E7FE4D65DB98F8BF56D255257EAD8B6E;
defparam prom_inst_0.INIT_RAM_10 = 256'h14E9F4E55386431BEE78E4EFA9F861BEE52677BB5510524EE4D55495CACA3B89;
defparam prom_inst_0.INIT_RAM_11 = 256'h65549BA9455C566F55C674924B509D527EED4249494A15F5227CE1834EE24E19;
defparam prom_inst_0.INIT_RAM_12 = 256'h75BA94559768ED4C9622AF6E75CBC66F8855571BBB7AEC6D6A9E475B79D571C5;
defparam prom_inst_0.INIT_RAM_13 = 256'h955F8694E72394A1D719ED624593581712B59E79A0519E5E20AE8CE1B39393B3;
defparam prom_inst_0.INIT_RAM_14 = 256'h2B541792B8F7C657653D6609576669DD2C955E1B5454541D7214D4104224A2C5;
defparam prom_inst_0.INIT_RAM_15 = 256'hAAB03B12296D57B5AA4C6562249E17A34510DD466995D2C6549E8D59669D093B;
defparam prom_inst_0.INIT_RAM_16 = 256'hA4770A9587CF722E755C55F5C65F16DB5476753B6D4EBBD59E9DDED45293DC67;
defparam prom_inst_0.INIT_RAM_17 = 256'h5852DCC2FDA3A74182363396162955DB29453B862422098D95D3995AB1577DD8;
defparam prom_inst_0.INIT_RAM_18 = 256'h98ED253B68924C7A31BED542792C3BC239277D450F3A8ED00B08B79D1282F9AE;
defparam prom_inst_0.INIT_RAM_19 = 256'h96F692AF552CA6E7ED25879E7B68A29F13D2F6B964B2B9FB4985A97F6908A2AA;
defparam prom_inst_0.INIT_RAM_1A = 256'h7B004B7B95DAEED6ABB4B8491BB46075B1997BDA4A57C62795DC7355EDDDE5CA;
defparam prom_inst_0.INIT_RAM_1B = 256'hEB68BA2E29421596B4964B3D7CF2B9165558A795C46DAF4535F5C575F95E5789;
defparam prom_inst_0.INIT_RAM_1C = 256'h3AAE25A9EA38958AA9D396254ADF69EE4D6D7557287DFF6F4ACE09ABEE4D5686;
defparam prom_inst_0.INIT_RAM_1D = 256'h8656E6965E5AFDDDD6D93D46A6557C978CA5B715575567597D46EA6BBEAAAA66;
defparam prom_inst_0.INIT_RAM_1E = 256'hA50F1A2DDF7956EFB94ACE75755F7E320BECAD58F63FA455B5D7DDB5579C2381;
defparam prom_inst_0.INIT_RAM_1F = 256'h18A0865257728C8B677657D9DC952BC6761B9E4F4577D47BFB5576BBF873FF6F;
defparam prom_inst_0.INIT_RAM_20 = 256'h757C65561525FBD1B52D64791555E25729D6574BFF3B80B93B57B5A65757914B;
defparam prom_inst_0.INIT_RAM_21 = 256'h15CDD08D71B5AF27CD8905727A9916B18EEEC8ED86D77B6595486567D38ACDF5;
defparam prom_inst_0.INIT_RAM_22 = 256'h218F52CEA797B2907795B5549154142D5FB9BBDE7BFF5E6BDAD4B78D29F9095C;
defparam prom_inst_0.INIT_RAM_23 = 256'h7959195D97155565E7B79EE5BBBB56561BCDD0F5F556EF713D5869857F0BF2C9;
defparam prom_inst_0.INIT_RAM_24 = 256'hA4657F52A22EAECBE4AD6FFD4615D765B985F9179955557D7922FD5E85319579;
defparam prom_inst_0.INIT_RAM_25 = 256'h7BEB75CAC14E414826975A95F4AAD77BD2CE5B9F31B984F79975E892B5F4A658;
defparam prom_inst_0.INIT_RAM_26 = 256'h344AF6EC15555447D744D52433BBE275EB5DAF5296B6D7F72D77B73E7FBAD75B;
defparam prom_inst_0.INIT_RAM_27 = 256'hCA549FAD52B44F1D667BFA13BBEDBDD1C71DA75F96958A56667B75967C4D4149;
defparam prom_inst_0.INIT_RAM_28 = 256'h2436C72526FE5D795122EF561490E27F26F7699A59AEF8855178AFF54528D7EE;
defparam prom_inst_0.INIT_RAM_29 = 256'h5A572513D14CD099755F745371D3990D18A7A5EEFD215CF6C294DD7D74F426E6;
defparam prom_inst_0.INIT_RAM_2A = 256'hC9465D7D7348DB48CD55F5BF6965D3D6D653AD7578BA56557CF4209D5E33574F;
defparam prom_inst_0.INIT_RAM_2B = 256'h02000DF4AE634412E452D05BDF954B6888D25B7F2CDBEBFB34E5648D2B5A54B5;
defparam prom_inst_0.INIT_RAM_2C = 256'hB55B69159510D16462F189291AD027F3FFBD1F69C9BA889D79F73FE55DBEBF93;
defparam prom_inst_0.INIT_RAM_2D = 256'h4B15D4107576D621F3FFBD79D4999F26EF955B574014B79E48C5584575641061;
defparam prom_inst_0.INIT_RAM_2E = 256'h7C99B2D83C917AC4FE545FB92B2BC7DFBFD6D15B52BAC8954AFFD3ACEB3AC39E;
defparam prom_inst_0.INIT_RAM_2F = 256'h957BBB9577916FD7779D6DCA74C53CB234412C50FE78D24C11674A8CC5349DF1;
defparam prom_inst_0.INIT_RAM_30 = 256'h58A45C3B5B098CB420389C53FF54BCAC9C8D7146747175CB1BFF7FFFF9D467F8;
defparam prom_inst_0.INIT_RAM_31 = 256'h7D14A18529034E0FCE1A56D54E63A9257FF473B8E5909092B70921015475C818;
defparam prom_inst_0.INIT_RAM_32 = 256'h185B5552CDC5DB5F4662D9E2C565A7D2F6D151F2BFF6D79D4F55D275574D5754;
defparam prom_inst_0.INIT_RAM_33 = 256'hDA6EDA278A58AD6565C7D7B52FE7EBECE71578A72E966955AC4892179D4111B5;
defparam prom_inst_0.INIT_RAM_34 = 256'h48165E71355356EC7955B4BAAE315E69D5F504200C318005E737D055FCEAEA38;
defparam prom_inst_0.INIT_RAM_35 = 256'hED59715B754040FFA8228AEC0827906DB757556176D72A237224A5B51D655857;
defparam prom_inst_0.INIT_RAM_36 = 256'hFF335D13CBA012B2F9F175FF51862E0697D7FF2E8279376271CD65F5955455B9;
defparam prom_inst_0.INIT_RAM_37 = 256'h5F75DE94F0D8AE7017E3F745DF747C51FBC55F5D5375A575F75D5DF45194933F;
defparam prom_inst_0.INIT_RAM_38 = 256'hB96D474F6D653B75B27503A232719190DB28F97D84155A5512992D20C63D75F5;
defparam prom_inst_0.INIT_RAM_39 = 256'hC4512441DCBA2BBFCCBA2BBBD97FF72084289F7208240A65B555BFB593D6D657;
defparam prom_inst_0.INIT_RAM_3A = 256'h2B545EE11D49A441EF65FFC7C8AFC02FC185996D557A545EDC8AE4A0922BCD55;
defparam prom_inst_0.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7E521154CA20C35FD5727A092;
defparam prom_inst_0.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[29:0],dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 2;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h0268C2F801D8C0C243000FC3880F092E1252FFFFFFFFFFFFFFC8FFC4FFCCFF20;
defparam prom_inst_1.INIT_RAM_01 = 256'hD1C012FBFFC3D1C3112C60C89C1C0C03008CA8E78C280AE262C1D1C0C200003F;
defparam prom_inst_1.INIT_RAM_02 = 256'h2F7E0106105CF210E4003104FFFFFF0E4308410C10C7CB2DC107048000AC0EFF;
defparam prom_inst_1.INIT_RAM_03 = 256'h8187C82CCBC2CC5BCCCBC39B3213C1970210D6E9C6330A37739C008677CB00C3;
defparam prom_inst_1.INIT_RAM_04 = 256'hFE775171E5FA98A6BB24226940D23DC2D730B2098221988CB1D050800A0B5105;
defparam prom_inst_1.INIT_RAM_05 = 256'h14450DBF964C1EF501B5B1561F7F5CD34C541353446D375744E54E116735D577;
defparam prom_inst_1.INIT_RAM_06 = 256'h377B256534C783097DC00C3910407B4FCDCFB851FD980DD815D404F01C4B7C78;
defparam prom_inst_1.INIT_RAM_07 = 256'hC9DB5DA99AEE62ACCBB3FAF1812EDEEE6A6AEA3F3EF6EC5B59855DE199200C51;
defparam prom_inst_1.INIT_RAM_08 = 256'h1000110F2234B5BDBAA09E849EA90234E4FC60B04CAF5C433D6350DF7174C7E7;
defparam prom_inst_1.INIT_RAM_09 = 256'h0C0390F894BFD37A13972A35C14D8A0C5E4A2244C33842100BB0E03043F00000;
defparam prom_inst_1.INIT_RAM_0A = 256'h9C0D6405B6356F9D64C0F0B623233977097F022DC5E75F97F548C87ECB0C30C7;
defparam prom_inst_1.INIT_RAM_0B = 256'h385F4C293D0900270F0164E2175106100006206D80A78088517022A5162479B5;
defparam prom_inst_1.INIT_RAM_0C = 256'h2FF43426948D48F11C0C05CD7F82500021F1088E0C30A9F2060208811C21C3BD;
defparam prom_inst_1.INIT_RAM_0D = 256'h29A7505010B7A7002A89416B523CA762EDA6194ADD512DD52D63F571114BDE3D;
defparam prom_inst_1.INIT_RAM_0E = 256'h68DE7ABE6F369E235CD64A4BF8C8C4442F5D85E585F6A75D25420D2A000460C1;
defparam prom_inst_1.INIT_RAM_0F = 256'hB7003BE56424668D401297260CE30D4B5D85D00271EE68D800B13F155034AD2F;
defparam prom_inst_1.INIT_RAM_10 = 256'h008BF0A5820E60A125F6CEC484F6CB875C3BE44EF638DA213275B08EC8CA3F7B;
defparam prom_inst_1.INIT_RAM_11 = 256'hCE7A0EF80144DCD6F7024396EE8805CE4399AC1B8032F48C071083A0223EC839;
defparam prom_inst_1.INIT_RAM_12 = 256'hA028086D8EA82AFCE632F25384875C7886649E024C9931C66BC08C440915174D;
defparam prom_inst_1.INIT_RAM_13 = 256'h39EEE3E0CB1398413A0069237298410232320212ADD08D00100F6638D0F8CADB;
defparam prom_inst_1.INIT_RAM_14 = 256'h417882949BCE1C9EBDDB2A199EBDA90A1C4AA8797A149C090B82F4002E33AE5F;
defparam prom_inst_1.INIT_RAM_15 = 256'h88CA9DA138324510A4700107F97D10FA865F05C26F8D1F0251B3A246D6601032;
defparam prom_inst_1.INIT_RAM_16 = 256'hFDEC3E3BAEA6EEF74E07D87C3C78F3B1712C173A45C24C1299B7C00DD095BEE4;
defparam prom_inst_1.INIT_RAM_17 = 256'hFC41B242A0373EDB4266518A4A12EBA109DCCAFAF72BC9EBA7ACAA7B97DE9BAA;
defparam prom_inst_1.INIT_RAM_18 = 256'h760BE05108B410F13538273C5737C0C2C9929B4DE3D370B6092BC17DB180D7B5;
defparam prom_inst_1.INIT_RAM_19 = 256'h7250B6359F2426A672607D7FC10B6FD3BDBF0034270DA99C987DCF66CBE0833C;
defparam prom_inst_1.INIT_RAM_1A = 256'h039034C0E78C931274CF1BCB53D806782705A242389E3CFDA787CAE7B1388FB6;
defparam prom_inst_1.INIT_RAM_1B = 256'h693F0FE11F5B8184EDB3469B7270977EE793F0A8080B24C0BD4C7C7D13536417;
defparam prom_inst_1.INIT_RAM_1C = 256'hABFAF48FE3FAE707C23A9279C0F4291325E1C1DC268CC428C2C7B48F06C2721E;
defparam prom_inst_1.INIT_RAM_1D = 256'hEF6938C7C3BC09390AB7DBCFA3A77461342227B8DDF46DF69BCF0539F2B28F2F;
defparam prom_inst_1.INIT_RAM_1E = 256'hED3B868844C35130CF40EE78DD0DB742976C2D22C8B3C3209D5E089F776AFADB;
defparam prom_inst_1.INIT_RAM_1F = 256'h1A700EC29F303C1748F69FCA3DA703DE8D035E36E9EC03FBE9F7DE54F43DCF20;
defparam prom_inst_1.INIT_RAM_20 = 256'hAD50260860C880021718C8306D24E114285F4408001862060972A3961170A103;
defparam prom_inst_1.INIT_RAM_21 = 256'h350002089080806F00B81103095B451080132C42C65E3AB3944C0049B2BF7920;
defparam prom_inst_1.INIT_RAM_22 = 256'h30BCCA8E3CF190A023A1A8A237223405D04C4F46002AAB29045C63134AA1030A;
defparam prom_inst_1.INIT_RAM_23 = 256'h1010727B31F4446460009D36884CDFB47000356E6F739A7B9B5B071CCD098100;
defparam prom_inst_1.INIT_RAM_24 = 256'h610FA09CC08E8E7CF41A000510780F4F4C1D0D60F2EBDF4FD4035B41C1C09800;
defparam prom_inst_1.INIT_RAM_25 = 256'h28031786884E402064474AC882025CB7CA8E4D10DFD7AF4CF2C43CC1177C0320;
defparam prom_inst_1.INIT_RAM_26 = 256'h6887A79A709500845C285CAD904C31441978A8A1C204664CE5E3A001D0C65E3A;
defparam prom_inst_1.INIT_RAM_27 = 256'h86822485CAE848F8ADC002BF4C3021302CB8643030B4BD4A7DCEC29408801F2B;
defparam prom_inst_1.INIT_RAM_28 = 256'hE56F90245C80C0F3F619104074C9AB735C801972CE930B934C9C072D32105EB9;
defparam prom_inst_1.INIT_RAM_29 = 256'hD69E3532133031178426E80ACBF71FBF51F419D30D64E263C1F5009B4F6D2BF6;
defparam prom_inst_1.INIT_RAM_2A = 256'h6B4B05E5EF60593A67C04DC4E0813DB67CCCA7A9EB1A3CE7436CC1139620C4F6;
defparam prom_inst_1.INIT_RAM_2B = 256'h13313538715D329453165E63E5A63340E6D6419C9FEC6CED351B379144DC214C;
defparam prom_inst_1.INIT_RAM_2C = 256'h61751B41F51101332E5729102600147BE7BEBF950C84A46EDBED3DF32EC6CCDC;
defparam prom_inst_1.INIT_RAM_2D = 256'h49705C0417B2214F7BE7BE28A39527B564C8561720032224CE5C0200BC7C002F;
defparam prom_inst_1.INIT_RAM_2E = 256'hA6B59152B4CCD6671C13170221296B65B656FE010210CCFD48DF83380E13953F;
defparam prom_inst_1.INIT_RAM_2F = 256'h4884C4C8A220893A4290AA4F205DC441330095ECDF2A4E704C7D78664DC504D7;
defparam prom_inst_1.INIT_RAM_30 = 256'h2AF328CA87C5774CB8DEB4D9DD8068E8E8E2BAEB22975C59AFF590F75C8A0419;
defparam prom_inst_1.INIT_RAM_31 = 256'hA7C28C7D92126EFCE46A9FB9E478BEA9FF55E9AE67EA30A92A0A388087D9A6FC;
defparam prom_inst_1.INIT_RAM_32 = 256'hC7E463246FE008DDF6E136415D3121B9E0B5193151670175EC02F11F55A5B1F6;
defparam prom_inst_1.INIT_RAM_33 = 256'hF60916219F98FA260C025C4E0AF878D9D1355BD41360644F3782E2C045EFDF8D;
defparam prom_inst_1.INIT_RAM_34 = 256'hFAC8083CBD09D604F65594992A9704E05E1C00204210400A81BC452010260977;
defparam prom_inst_1.INIT_RAM_35 = 256'h35C6D355170000FFE8E1A37C5C98802BA1F6D0137D452119D0B39BA085DB06D5;
defparam prom_inst_1.INIT_RAM_36 = 256'h65C31FDD9274C161FE937ED6032311CE6D3B5115631332E317907D4C6D56C053;
defparam prom_inst_1.INIT_RAM_37 = 256'h09D72E5C466576700BAC81D1FB1D55DF915D7B1B09D76C17E085DFA2422A4A86;
defparam prom_inst_1.INIT_RAM_38 = 256'hC4678CC8E7CE124F4F9803AFE73BB787CE729AA8BF4546E00E8CE7EB5D88D797;
defparam prom_inst_1.INIT_RAM_39 = 256'hEEDBAEC0A454AF7FEC54AF520C11C008E43B38008ECF8E319F78009F3DB67CCC;
defparam prom_inst_1.INIT_RAM_3A = 256'h3883DA93FD87AFC0883047044CC89908A8E44C67DD0783DAACEB56B87A382DAA;
defparam prom_inst_1.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC5E3817200300803CD0BB38FE;
defparam prom_inst_1.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[29:0],dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 2;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hA2B8E32F85CFE3E3FBA22FEBA72F8F1A21B1FFFFFFFFFFFFFFC8FFCCFFC4FF33;
defparam prom_inst_2.INIT_RAM_01 = 256'h29C48DC30C23630C299E3302D85E3A2BA2EA360F0E307E01CBC5CCE3E38B88BF;
defparam prom_inst_2.INIT_RAM_02 = 256'hCC23306D8A095389C0809304FFFFFF2E6E8AFBEBBBAA8002BA6EB2C81BD040C3;
defparam prom_inst_2.INIT_RAM_03 = 256'hC8022B50E72502A79ED7998099BB1040A603F1E8CC8304FE333EA88C40140AFA;
defparam prom_inst_2.INIT_RAM_04 = 256'h65656649774755455746584773BBEA003AEE8BAFFA2BABF80BBB9810BD00AEBB;
defparam prom_inst_2.INIT_RAM_05 = 256'h5114510010504000440004041040511411511404510144100101501050400767;
defparam prom_inst_2.INIT_RAM_06 = 256'h4040400044041414001551404550401FD006A915001850181404400100504041;
defparam prom_inst_2.INIT_RAM_07 = 256'h14DF5D76C088040665595891D5C45848048C0808CC8C44809019020242404065;
defparam prom_inst_2.INIT_RAM_08 = 256'h0000110701017D4E545544767743003078784110C0401054410E041040011000;
defparam prom_inst_2.INIT_RAM_09 = 256'h06A88416E35F97B009A02030082080800202FAA203BC22AC0082A8EF2BFA0000;
defparam prom_inst_2.INIT_RAM_0A = 256'h12784DD0448C4F10502AF9418C8E373B200F6A5021041344F423232141245045;
defparam prom_inst_2.INIT_RAM_0B = 256'hBA02AE8BB0A84EE12EA84EEA84036DA6EE9E9A020A60366A100419A24C0F048F;
defparam prom_inst_2.INIT_RAM_0C = 256'h87F23EF0302C22FA42FA412C4F262AA79AABAEE6269A6228AE9AAA6BBAA0873A;
defparam prom_inst_2.INIT_RAM_0D = 256'h8C0F085BCC32345938B088CD85BE8400F07D688CEC2FA3627C9BF0100527C1FC;
defparam prom_inst_2.INIT_RAM_0E = 256'h30CC730CCC320F8E10C8E313C02382A00C100120013323100088CF8C556A3118;
defparam prom_inst_2.INIT_RAM_0F = 256'h143BF330C2F2336F3538F304AEC71CC310010A7F34CF06C0194A983908730CC7;
defparam prom_inst_2.INIT_RAM_10 = 256'hE626F62628A2801F5138003D4134F12F12B72A64C00300F888808020A3A30F94;
defparam prom_inst_2.INIT_RAM_11 = 256'h00400EF50127202000AAA8A102D32022A9990048C28888027B32288C8435228A;
defparam prom_inst_2.INIT_RAM_12 = 256'h2AA05A222232A8FFC4B7FA080A800DB0444512AA6623B8CCCFE603029AF49872;
defparam prom_inst_2.INIT_RAM_13 = 256'h010DD3CA2008A23182AA6849F98030ACC8E9A698CEFA8FA6327FD231D1C8D9D1;
defparam prom_inst_2.INIT_RAM_14 = 256'h340089A3575E8C12318088BA1230422917799A3405B9101841194814117AC760;
defparam prom_inst_2.INIT_RAM_15 = 256'h32E33C300CB86039C8FAA8413C8D0416A249A02A8820F3AAA04020410412BA9A;
defparam prom_inst_2.INIT_RAM_16 = 256'hF1082C83308008336097227271C9C70408814098102A66AAA10066B13BDC030C;
defparam prom_inst_2.INIT_RAM_17 = 256'h0EA330EF125250DF2F0808EAEAB51023BE1013C4B8CB32C3048C244218028000;
defparam prom_inst_2.INIT_RAM_18 = 256'h001418339C0FBEAEAA72048004B314AF029E806302244537BC8C0C4B38EF8431;
defparam prom_inst_2.INIT_RAM_19 = 256'h4079C0B1104EF482F891004F139C8BD8C80329EEA8CB20BE2402D4B0141233BD;
defparam prom_inst_2.INIT_RAM_1A = 256'h98C04810C4A299841EE23200AEAABF32502D32E74C1288B204A72604118694A3;
defparam prom_inst_2.INIT_RAM_1B = 256'h79304C1D1C1FC9A60040468002CBFC430412F9B12AA8C71252727242987B7008;
defparam prom_inst_2.INIT_RAM_1C = 256'h62C0B1054360C46B34C644912F84888855002002774A414FEF53662CCF30488D;
defparam prom_inst_2.INIT_RAM_1D = 256'hCB6A80049843298AAA8080109FC400098EFAA8C2010A613480101D72C4B52C8B;
defparam prom_inst_2.INIT_RAM_1E = 256'hC57E473E7718C48AD46F94820347C0C7E576F0AF3AC887B303628B000EC8B2D2;
defparam prom_inst_2.INIT_RAM_1F = 256'h7274D4E7100BF32453051024C144BC8D30BEC2200122072CB000115C720D8CC2;
defparam prom_inst_2.INIT_RAM_20 = 256'h305AE8AA1AB2AED5003A6A9A020A600A6100D694AA6276277009A998A40A969E;
defparam prom_inst_2.INIT_RAM_21 = 256'h4BBB0740DBEE2A10BB1304457160303BD899BDCBD4029A79B946EA68072F7AAC;
defparam prom_inst_2.INIT_RAM_22 = 256'h1471E2A651473BF0A989A0A703D549503A666C15EEEA29891400E988358373E9;
defparam prom_inst_2.INIT_RAM_23 = 256'hAAAA304809C6AAAAAAAAAAB03E660045453B830200099A8C80421051C8BDC4EE;
defparam prom_inst_2.INIT_RAM_24 = 256'hE850EA12D8D8D8CEC988BBAE89C152902272AC71451000030E7380114BEAA2AA;
defparam prom_inst_2.INIT_RAM_25 = 256'h990600AEAEA6828AE1CF1173A8950230A2A6F36000C40571452114EB8072F3AA;
defparam prom_inst_2.INIT_RAM_26 = 256'h250AA888F906F1AA029A02203E66B31C500A2A002897CB718029A1043AD4029A;
defparam prom_inst_2.INIT_RAM_27 = 256'hAE2881C0221549CAA014442A22BA728A410A2989850154AAB0202AA18ABB8088;
defparam prom_inst_2.INIT_RAM_28 = 256'h4053905551C61524000A8AA1C01D1F8A51C389840C59A114103EF65040B80288;
defparam prom_inst_2.INIT_RAM_29 = 256'h10121D48144208D80120238605442C5842F2C6ABA505013710F10B8062014BD0;
defparam prom_inst_2.INIT_RAM_2A = 256'h90D746252E7563ACF41271471A15880400104031213C0004620238D810A80620;
defparam prom_inst_2.INIT_RAM_2B = 256'h30011608B87FAB11CA98C74C35E0AE72C7A453CA911E5E5C661C20399417AB63;
defparam prom_inst_2.INIT_RAM_2C = 256'h49449C1141F4D33A86D8383B16001C1D75C72A0601474401D75C6BBA80E4E4C0;
defparam prom_inst_2.INIT_RAM_2D = 256'h018460121405090E1D75C4BE9BA579298EEAA7A6940BABF608612D4C53501018;
defparam prom_inst_2.INIT_RAM_2E = 256'h2D06304F90AAD0F014BAA53F9D9C7875D75B7F87F9DDC60CA75288FA7E9FBD8E;
defparam prom_inst_2.INIT_RAM_2F = 256'h2922266A2AAAA9C2AAAAA8CBAB6184E0CA81060C5BACEB00EA50040F7004EE98;
defparam prom_inst_2.INIT_RAM_30 = 256'hADFA80ED2441D76177E90723502878F8F8F8973EA8D89A63C91CFA7DCEA10274;
defparam prom_inst_2.INIT_RAM_31 = 256'h24358F637D379C05985910C118362D110944272DCEC535466A5673C2361FDD0D;
defparam prom_inst_2.INIT_RAM_32 = 256'hF618D0D2D4350539390FAD7B62AA59C4A941A51D003511C51C494DD060353D0C;
defparam prom_inst_2.INIT_RAM_33 = 256'hAD3B8D4DCB63F9C1C0BA62411A1E5E5C89C61CB2FADC19EF3364DBCC0610D053;
defparam prom_inst_2.INIT_RAM_34 = 256'h076AAA9E534705F73F143035D0D8461A5292000082242009EB52D70BBBB11123;
defparam prom_inst_2.INIT_RAM_35 = 256'hB5251C95540000FFE9EAC2E3D814005C490534D4412D1007113AD4B4C5144505;
defparam prom_inst_2.INIT_RAM_36 = 256'hEDCB9853727E632309DC400129C302E751C00B020998B9F99842527252C4D318;
defparam prom_inst_2.INIT_RAM_37 = 256'h851401262D1A17300058691D0593F6104F614594471471181405105AD666394E;
defparam prom_inst_2.INIT_RAM_38 = 256'hE24021A180008F61431003AB3B73737F8F23D01661E96714064EB4DF61C51894;
defparam prom_inst_2.INIT_RAM_39 = 256'h740594028300CC803300CC862A3BAECBF23D4EECBF508FA80002EE000804001C;
defparam prom_inst_2.INIT_RAM_3A = 256'hB52723BDCBB5170298A8EEE2C3D107D108F12A00004927238DD3133750B5DBAA;
defparam prom_inst_2.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCC103CB2227300023E4493F7DC;
defparam prom_inst_2.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[29:0],dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 2;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h04F0C47FEF00C40470000340030313B03BF0FFFFFFFFFFFFFFCBFFC7FFCBFF2F;
defparam prom_inst_3.INIT_RAM_01 = 256'hF1C71130C307F1CB001C42C0DEE0484000CCF0F9CC4EFC7BFF6E00C40413000D;
defparam prom_inst_3.INIT_RAM_02 = 256'h0F0F1C0411002F10407033C7FFFFFF0045105545514550015545545150107C30;
defparam prom_inst_3.INIT_RAM_03 = 256'h5070C82CC0F2C0D96403C2032033C2CF202D970CF832CB6452E420B871CB1003;
defparam prom_inst_3.INIT_RAM_04 = 256'h0200200210032221002311312151554015555140004155550401515501005515;
defparam prom_inst_3.INIT_RAM_05 = 256'hD575D55755D755D55D5D5D7575775D5D755755D55775D5D7575D5757575D7110;
defparam prom_inst_3.INIT_RAM_06 = 256'hD755D5D5D75D75D75D75D75D75D75D7A9D7EA95D7571777175D5755D57575755;
defparam prom_inst_3.INIT_RAM_07 = 256'h114D245040CC40C8888444C808CC4C8CC844880884C48A1715715C5C5C5D75C5;
defparam prom_inst_3.INIT_RAM_08 = 256'hC7000003339D87B9A0AD9CA890B40304D4D4F30CF55555555550555555555504;
defparam prom_inst_3.INIT_RAM_09 = 256'h0080030F13EC6CC00033C313FF3CB3C03F3F95C47B1001550050505540F20C30;
defparam prom_inst_3.INIT_RAM_0A = 256'h1C0BC3F47C3C701C71C8F0B20F22C0C91CFF082C83C73D0F0403C80C00000000;
defparam prom_inst_3.INIT_RAM_0B = 256'h153D44321520F473CA007857033E04204437033F3C03FC052CF00032F8FF2CFE;
defparam prom_inst_3.INIT_RAM_0C = 256'hF833D8C0E0CD3CD200C8B3C0F0C0F00001630CC8C00001E00C002001188CFCC5;
defparam prom_inst_3.INIT_RAM_0D = 256'hF83947730F73CC03DFF4BCB9CF74073ED4F83CBB742E3572DCB75333233CCB34;
defparam prom_inst_3.INIT_RAM_0E = 256'h0DC333CF0F32CD223C07880DD0C88081CF3C73C073D0C03C7032022300083C00;
defparam prom_inst_3.INIT_RAM_0F = 256'hCBF303E0F0C483CFF3E233C7CB79E4B03C73C0052C1D1CC7FCB20B0FCB30CC37;
defparam prom_inst_3.INIT_RAM_10 = 256'hFC87F08FF208C71E03DC7078085C30C93F00FC44FCB1C7911C7CFF0F8808CDC7;
defparam prom_inst_3.INIT_RAM_11 = 256'h3C70C2D583F3F3E3CFC8F033C3F2F3C0C1130FCB0000FF0C043C8207CB31C823;
defparam prom_inst_3.INIT_RAM_12 = 256'hF003F53F0F1C8F00C73CD3D108C10F30EFC01F23442E10F833402CE3033FCB3F;
defparam prom_inst_3.INIT_RAM_13 = 256'hF1F1F77C81023C8C3F200C3090070C8CF2200000B2723F00FC8CC03CFCC0C0FF;
defparam prom_inst_3.INIT_RAM_14 = 256'h3CF00033D967CF1C3F0FC7331C3C30FC04F0053CF23F1C0030DC3C0A07B0032C;
defparam prom_inst_3.INIT_RAM_15 = 256'h3CCEE55000CC01E00F908C30BCBCC30C53CF33C8CF0F38C8FCF02C00C30F3323;
defparam prom_inst_3.INIT_RAM_16 = 256'hD3C7CC30D123C7B50FF3FF3F3C3CFC1CF007CF2073C8443031CF00F3F338F2CF;
defparam prom_inst_3.INIT_RAM_17 = 256'hC0803F8C2F2E2CF88C0F12000001C73E333F1CC33C3B0EF3C7032C73CB3C8F2E;
defparam prom_inst_3.INIT_RAM_18 = 256'h31CB133E000554551542C7C70F041E0C1FBC0F0F1C0CC73E31203CFBC20C8F03;
defparam prom_inst_3.INIT_RAM_19 = 256'h036003351C38CCFC90BF1CF01E00F37CB0F2F02C0CB03F242F1F0BC3C72C8034;
defparam prom_inst_3.INIT_RAM_1A = 256'h00B00F1EC7C0D1030841E3C05554554F2C4B1F80CB1CC730C733F2C70FC0C700;
defparam prom_inst_3.INIT_RAM_1B = 256'h6830CC3B04F770001CF0C00F0FA30CF1C70CD030D48CB3EF0F3F3F1FCFF1F0CB;
defparam prom_inst_3.INIT_RAM_1C = 256'h2CC7B0C0773DC7032CF2C301CC8F031153D7333CE50C60B60C73EC04393C700F;
defparam prom_inst_3.INIT_RAM_1D = 256'hFB35104C8CB3FC3FC0CF0F3CF347D03CF8C03CBF3CFC03D30F3CFB2ECBB1CCBB;
defparam prom_inst_3.INIT_RAM_1E = 256'h80CACDE773CFFD104FCC83C83FF2443E5110C1396E58311F0F3FFF0CFEF3BCCC;
defparam prom_inst_3.INIT_RAM_1F = 256'h1CD0CB001D8303CCF3CF1D3CF3C7318F3D32F203F1C3F1C510CF3D0BBEE0B070;
defparam prom_inst_3.INIT_RAM_20 = 256'h3FDCCFC0200FC471CF0005033FCC003F1F3C8FC3001C90C90CF0300F00F01702;
defparam prom_inst_3.INIT_RAM_21 = 256'hBF1133C04304003D110F00300E3D70E30B1124B24F3F03003CC0CC00F1CD4FFF;
defparam prom_inst_3.INIT_RAM_22 = 256'h059640C83CF1E30030303300D4CCBCF3FC470547C4430D01033C000F3CD73CFC;
defparam prom_inst_3.INIT_RAM_23 = 256'h03033C70FCFC0C0C00303510E4473CBC31D1D63C3CFD13CB0FF3030C7930B84C;
defparam prom_inst_3.INIT_RAM_24 = 256'hC007731CC7878784CD03D10700BF3DC7472F0700F1C73CF2D8088F0C3E423F03;
defparam prom_inst_3.INIT_RAM_25 = 256'h00730FCCCCC8C000CC8E0C3FC00F3C3100C8F22C0CCF303CF1C0C3730F3CC000;
defparam prom_inst_3.INIT_RAM_26 = 256'h45010D139FFFFF5F3FF53C05EC441BC00CFC0C0070038D3C73F03C31E0433F03;
defparam prom_inst_3.INIT_RAM_27 = 256'h0CF004F3C045FCFC03CF00C1441F1FCC3CFC0CFCFC70C2C0D3F1F03CF151CF01;
defparam prom_inst_3.INIT_RAM_28 = 256'h303DC78F3C73F3D1D40510FCBC0479DE3C7D0031C31100C3C8E4C63F23333C11;
defparam prom_inst_3.INIT_RAM_29 = 256'hC31C0C31C32CB203DFC3FDF2C073CC0F3CDF535104F0F769708C4F0F0C3CB3CC;
defparam prom_inst_3.INIT_RAM_2A = 256'h43F3F3F3F01E3E0393FC3C73C0CC30FC33CB03D1C0E433C70C3C4203C3A2F0C3;
defparam prom_inst_3.INIT_RAM_2B = 256'hC8CCC3DAD13E01CF600F953D9443022FCD553E5943646465A3C300C0F0CB020F;
defparam prom_inst_3.INIT_RAM_2C = 256'h10710F3C7F78C810038B8993862003451451C930C150CC365965991036464643;
defparam prom_inst_3.INIT_RAM_2D = 256'h0CBF3C080FD57CF445145203C033D40CF840F23214003011C32FC4200F1C0A0F;
defparam prom_inst_3.INIT_RAM_2E = 256'hC433DB2D86804B90C3C030E910111114510F01FCF1030C77C456D1104411007C;
defparam prom_inst_3.INIT_RAM_2F = 256'h00C44440F0140CFFF03C0F6D032CB200500082F38303800F001D0CF93C33FB0B;
defparam prom_inst_3.INIT_RAM_30 = 256'h02D03324F0C0F10E81D833FE55FF9393939380F6034BC82E78405004040C3010;
defparam prom_inst_3.INIT_RAM_31 = 256'hF3FCF33F3C39CB068F031CF1CF73CC31D153C2CCBCF2C3C2F33C0E40F2C76077;
defparam prom_inst_3.INIT_RAM_32 = 256'h33C7C3CB837240F8FC3000702F0320B8BCB233D38811FCB3CBFC33CBFD97CCBF;
defparam prom_inst_3.INIT_RAM_33 = 256'h0030103CF33CD0F0B31F3C0CF06464640CFFCF00000B00F0042CCB2C03C7070F;
defparam prom_inst_3.INIT_RAM_34 = 256'hF0C0C0C70FF1FC73DDF3E0E1CB4BF3C03FCC00004300A80C7E0CC93D110C3300;
defparam prom_inst_3.INIT_RAM_35 = 256'h13F2CFF20F80A05F694B6145610B700F30F1FFCB1C4CB3B1CBB00B8203CBF1FC;
defparam prom_inst_3.INIT_RAM_36 = 256'h44F10B011ED048485D4F1C68812303042CF1A103B10F10710B0F1F3F2FFF3F0F;
defparam prom_inst_3.INIT_RAM_37 = 256'hF2CF93A781A18E1024CF30FC730FE2C73C2C7307F1CF3FCF3243C73171B96474;
defparam prom_inst_3.INIT_RAM_38 = 256'h47C3C9C9C33F210CB0FE01A56D9D49853D9134CC3C0C43D600EC03C32CF2CFCF;
defparam prom_inst_3.INIT_RAM_39 = 256'h00C030C0F4CC0CC014CC0CD0C0D18440D034F4440D3C0D030CFF470CF0FC33C7;
defparam prom_inst_3.INIT_RAM_3A = 256'h30F1F5F0760CB1C0C30346C04C0CC30CC0D000C33C30F1F5F0F3303CC330C600;
defparam prom_inst_3.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF3F0BB71C800C31FCC30C3CC7;
defparam prom_inst_3.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

endmodule //ROM8kB
